`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:43:24 04/20/2015 
// Design Name: 
// Module Name:    Principal 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Principal(
    input SW0,
    input BTN0,
    input V,
    output A,
    output B
    );
wire w1, w2, w3, w4, w5, w6
JK jk1()
nor (w1, SWO, w4, )

endmodule
